module sit
